module trnsfrm2d

// TEST
