module transform_2d
