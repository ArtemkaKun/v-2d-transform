module trnsfrm2d
